//edit2
module multi
(
    input [3:0] a,b,
  output reg [4:0] multi,
    input clk
  );
  
  
  always@(posedge clk)
    begin
      sum <= a * b;
    end
   
   
endmodule
