//edit2
module multi
(
    input [3:0] a,b,
    output reg [4:0] opp,
   // input clk
  );
  
  
  //always@(posedge clk)
   // begin
      opp <= a * b;
   // end
   
   
endmodule
