//edit2
